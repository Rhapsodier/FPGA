// ============================================================================
// BCD码转7段显示码
// ============================================================================
// 功能：将BCD码（0-9）转换为7段显示码
// 数码管类型：共阳极（0表示点亮，1表示熄灭）
// 段码顺序：seg7[6:0] = {g, f, e, d, c, b, a}
// 段位置：a为最顶端，顺时针依次为 b, c, d, e, f，g为中间横
// 实现：使用查找表（case语句）
// ============================================================================
module bcd_to_seg7 (
    input wire [3:0] bcd,
    output reg [6:0] seg7  // {g, f, e, d, c, b, a}
);

    always @(*) begin
        case (bcd)
            4'd0: seg7 = 7'b1000000;  // 0: 点亮 a,b,c,d,e,f，熄灭 g
            4'd1: seg7 = 7'b1111001;  // 1: 点亮 b,c，熄灭 a,d,e,f,g
            4'd2: seg7 = 7'b0100100;  // 2: 点亮 a,b,d,e,g，熄灭 c,f
            4'd3: seg7 = 7'b0110000;  // 3: 点亮 a,b,c,d,g，熄灭 e,f
            4'd4: seg7 = 7'b0011001;  // 4: 点亮 b,c,f,g，熄灭 a,d,e
            4'd5: seg7 = 7'b0010010;  // 5: 点亮 a,c,d,f,g，熄灭 b,e
            4'd6: seg7 = 7'b0000010;  // 6: 点亮 a,c,d,e,f,g，熄灭 b
            4'd7: seg7 = 7'b1111000;  // 7: 点亮 a,b,c，熄灭 d,e,f,g
            4'd8: seg7 = 7'b0000000;  // 8: 点亮 a,b,c,d,e,f,g
            4'd9: seg7 = 7'b0010000;  // 9: 点亮 a,b,c,d,f,g，熄灭 e
            default: seg7 = 7'b1111111;  // 其他：全灭
        endcase
    end

endmodule

